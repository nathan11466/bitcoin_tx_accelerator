// test bench for an accelerator

module accel_tb ();

  // accelerator outputs
  logic hash_done;
  logic mem_acc_read_en;
  logic mem_acc_write_en;
  logic [15:0] mem_acc_write_addr;
  logic [15:0] mem_acc_read_addr;
  logic [31:0] mem_acc_write_data;
  logic [255:0] hash;

  // accelerator inputs
  logic mem_listen_en;
  logic mem_acc_write_done;
  logic mem_acc_read_data_valid;
  logic [15:0] mem_listen_addr;
  logic [31:0] mem_listen_data;
  logic [511:0] mem_acc_read_data;
  logic clk, rst_n;

  // file handlers
  // f1: stores randomly generated block headers
  // f2: stores the SHA-256 hashes (generated by the accelerator)
  //     of the headers in f1
  integer f1, f2;

  // block header
  logic [511:0] temp_0; // applied at stage 1
  logic [511:0] temp_1; // applied at stage 2

  // Instantiate the accelerator
  accel accel0 (.hash_done(hash_done), .hash(hash), // output
                .mem_acc_read_addr(mem_acc_read_addr),
                .mem_acc_read_en(mem_acc_read_en),
                .mem_acc_write_en(mem_acc_write_en),
                .mem_acc_write_data(mem_acc_write_data),
                .mem_acc_write_addr(mem_acc_write_addr),
                .mem_listen_addr(mem_listen_addr), // input
                .mem_listen_en(mem_listen_en),
                .mem_listen_data(mem_listen_data),
                .mem_acc_read_data(mem_acc_read_data),
                .mem_acc_read_data_valid(mem_acc_read_data_valid),
                .mem_acc_write_done(mem_acc_write_done),
                .clk(clk), .rst_n(rst_n)
               );

  // Generate random block headers
  function automatic void generate_random_block_header(ref logic [511:0] header);
    header = {319'b0, 64'b10_1000_0000, 32'h{rand(), rand(), rand(), rand()}};
  endfunction

  // Write the hash value to the output file
  function void write_hash_to_file(integer file_handle, logic [255:0] hash);
    $fwrite(file_handle, "%h\n", hash);
  endfunction

  // Write the raw block header to the input file
  function void write_raw_block_header_to_file(integer file_handle, logic [511:0] header);
    $fwrite(file_handle, "%h\n", header);
  endfunction

  // Write the final hash value to the output file
  function void write_final_hash_to_file(integer file_handle, logic [255:0] hash);
    $fwrite(file_handle, "final hash = %h\n", hash);
  endfunction

  // Clock
  initial clk = 0;
  always #5 clk = ~clk;

  // Testing
  initial begin
    // Open the input and output files
    f1 = $fopen("hash_in.txt", "w");
    if (f1 == 0) begin
      $display("Error: Could not open input file");
      $stop;
    end
    f2 = $fopen("simu_out_accel.txt", "w");
    if (f2 == 0) begin
      $display("Error: Could not open output file");
      $stop;
    end

    // Reset
    rst_n = 0;
    mem_listen_en = 0;
    mem_acc_write_done = 0;
    mem_acc_read_data_valid = 0;
    mem_listen_addr = 0;
    mem_listen_data = 0;
    mem_acc_read_data = 0;

    @(negedge clk);
    rst_n = 1;
    @(posedge clk);

    for (int k = 0; k < 1000; k++) begin

      // Generate a random block header
      generate_random_block_header(temp_0);

      // Write the raw block header to the input file
      write_raw_block_header_to_file(f1, temp_0);
      $display("raw block header = %h\n", temp_0);

      // Stage 1
      // Start hashing
      mem_listen_en = 1;
      mem_listen_addr = 16'h5000;
      mem_listen_data = 32'b1;

      // Read the message from memory
      @(posedge clk); // @ READ_MSG_1
      mem_listen_en = 0;
      assert (mem_acc_read_en == 1)
      else   $error("error: mem_acc_read_en");
      assert (mem_acc_read_addr == 16'h1000)
      else   $error("error: mem_acc_read_addr");

      //
